LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY memoria IS
	PORT(
		entrada: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		saida: OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
END memoria;

ARCHITECTURE circ1 OF memoria IS
BEGIN
	WITH entrada SELECT
		saida <=	"00100000" WHEN "00000000",
					"10000111" WHEN "00000001",
					"00010000" WHEN "00000010",
					"10000010" WHEN "00000011",
					"00100000" WHEN "00000100",
					"10000000" WHEN "00000101",
					"10100000" WHEN "00000110",
					"01001010" WHEN "00000111",
					"00100000" WHEN "00001000",
					"10000001" WHEN "00001001",
					"10100000" WHEN "00001010",
					"01001010" WHEN "00001011",
					"01100000" WHEN "00001100",
					"00110000" WHEN "00001101",
					"10000110" WHEN "00001110",
					"00110000" WHEN "00001111",
					"10000000" WHEN "00010000",
					"10100000" WHEN "00010001",
					"01000110" WHEN "00010010",
					"10010000" WHEN "00010011",
					"00011111" WHEN "00010100",
					"00100000" WHEN "00010101",
					"10000000" WHEN "00010110",
					"00010000" WHEN "00010111",
					"10000011" WHEN "00011000",
					"00100000" WHEN "00011001",
					"10000001" WHEN "00011010",
					"00010000" WHEN "00011011",
					"10000100" WHEN "00011100",
					"10000000" WHEN "00011101",
					"00100111" WHEN "00011110",
					"00100000" WHEN "00011111",
					"10000001" WHEN "00100000",
					"00010000" WHEN "00100001",
					"10000011" WHEN "00100010",
					"00100000" WHEN "00100011",
					"10000000" WHEN "00100100",
					"00010000" WHEN "00100101",
					"10000100" WHEN "00100110",
					"00100000" WHEN "00100111",
					"10000011" WHEN "00101000",
					"00010000" WHEN "00101001",
					"10000010" WHEN "00101010",
					"00100000" WHEN "00101011",
					"10000010" WHEN "00101100",
					"00010000" WHEN "00101101",
					"10000101" WHEN "00101110",
					"00100000" WHEN "00101111",
					"10000100" WHEN "00110000",
					"01100000" WHEN "00110001",
					"00110000" WHEN "00110010",
					"10000110" WHEN "00110011",
					"00110000" WHEN "00110100",
					"10000101" WHEN "00110101",
					"00010000" WHEN "00110110",
					"10000101" WHEN "00110111",
					"10010000" WHEN "00111000",
					"00111110" WHEN "00111001",
					"10100000" WHEN "00111010",
					"01001010" WHEN "00111011",
					"10000000" WHEN "00111100",
					"00101111" WHEN "00111101",
					"00100000" WHEN "00111110",
					"10000010" WHEN "00111111",
					"00110000" WHEN "01000000",
					"10000011" WHEN "01000001",
					"00010000" WHEN "01000010",
					"10000010" WHEN "01000011",
					"10000000" WHEN "01000100",
					"00101011" WHEN "01000101",
					"00100000" WHEN "01000110",
					"10000000" WHEN "01000111",
					"00010000" WHEN "01001000",
					"10000010" WHEN "01001001",
					"11110000" WHEN "01001010",
					"00011110" WHEN "10000000",
					"00011110" WHEN "10000001",
					"00011110" WHEN "10000010",
					"00010100" WHEN "10000011",
					"00001111" WHEN "10000100",
					"00000001" WHEN "10000110",
					
					"00000000" WHEN OTHERS;
END circ1;