library verilog;
use verilog.vl_types.all;
entity final_work_vlg_vec_tst is
end final_work_vlg_vec_tst;
